`timescale 1ns / 1ns

// registers are 32 bits in RV32
`define REG_SIZE 31:0

// RV opcodes are 7 bits
`define OPCODE_SIZE 6:0

`include "../hw2a/divider_unsigned.sv"
`include "../hw2b/cla.sv"

module RegFile (
    input logic [4:0] rd,
    input logic [`REG_SIZE] rd_data,
    input logic [4:0] rs1,
    output logic [`REG_SIZE] rs1_data,
    input logic [4:0] rs2,
    output logic [`REG_SIZE] rs2_data,

    input logic clk,
    input logic we,
    input logic rst
);
  localparam int NumRegs = 32;
  logic [`REG_SIZE] reg_outs[NumRegs];

  // TODO: your code here

endmodule

module DatapathSingleCycle (
    input wire clk,
    input wire rst,
    output logic [`REG_SIZE] pc,
    input wire [`REG_SIZE] insn,
    // addr1 is a read-write port
    output wire [`REG_SIZE] addr1,
    input logic [`REG_SIZE] dout1,
    output wire [`REG_SIZE] din1,
    output wire [3:0] we1,
    output logic halt
);

  // components of the instruction
  wire [6:0] insn_funct7;
  wire [4:0] insn_rs2;
  wire [4:0] insn_rs1;
  wire [2:0] insn_funct3;
  wire [4:0] insn_rd;
  wire [`OPCODE_SIZE] insn_opcode;

  // split R-type instruction - see section 2.2 of RiscV spec
  assign {insn_funct7, insn_rs2, insn_rs1, insn_funct3, insn_rd, insn_opcode} = insn;

  // setup for I, S, B & J type instructions
  // I - short immediates and loads
  wire [11:0] imm_i;
  assign imm_i = insn[31:20];
  wire [ 4:0] imm_shamt = insn[24:20];

  // S - stores
  wire [11:0] imm_s;
  assign imm_s[11:5] = insn_funct7, imm_s[4:0] = insn_rd;

  // B - conditionals
  wire [12:0] imm_b;
  assign {imm_b[12], imm_b[10:5]} = insn_funct7, {imm_b[4:1], imm_b[11]} = insn_rd, imm_b[0] = 1'b0;

  // J - unconditional jumps
  wire [20:0] imm_j;
  assign {imm_j[20], imm_j[10:1], imm_j[11], imm_j[19:12], imm_j[0]} = {insn[31:12], 1'b0};

  wire [`REG_SIZE] imm_i_sext = {{20{imm_i[11]}}, imm_i[11:0]};
  wire [`REG_SIZE] imm_s_sext = {{20{imm_s[11]}}, imm_s[11:0]};
  wire [`REG_SIZE] imm_b_sext = {{19{imm_b[12]}}, imm_b[12:0]};
  wire [`REG_SIZE] imm_j_sext = {{11{imm_j[20]}}, imm_j[20:0]};

  // opcodes - see section 19 of RiscV spec
  localparam bit [`OPCODE_SIZE] OpLoad = 7'b00_000_11;
  localparam bit [`OPCODE_SIZE] OpStore = 7'b01_000_11;
  localparam bit [`OPCODE_SIZE] OpBranch = 7'b11_000_11;
  localparam bit [`OPCODE_SIZE] OpJalr = 7'b11_001_11;
  localparam bit [`OPCODE_SIZE] OpMiscMem = 7'b00_011_11;
  localparam bit [`OPCODE_SIZE] OpJal = 7'b11_011_11;

  localparam bit [`OPCODE_SIZE] OpRegImm = 7'b00_100_11;
  localparam bit [`OPCODE_SIZE] OpRegReg = 7'b01_100_11;
  localparam bit [`OPCODE_SIZE] OpEnviron = 7'b11_100_11;

  localparam bit [`OPCODE_SIZE] OpAuipc = 7'b00_101_11;
  localparam bit [`OPCODE_SIZE] OpLui = 7'b01_101_11;

  wire insn_lui = insn_opcode == OpLui;
  wire insn_auipc = insn_opcode == OpAuipc;
  wire insn_jal = insn_opcode == OpJal;
  wire insn_jalr = insn_opcode == OpJalr;

  wire insn_beq = insn_opcode == OpBranch && insn[14:12] == 3'b000;
  wire insn_bne = insn_opcode == OpBranch && insn[14:12] == 3'b001;
  wire insn_blt = insn_opcode == OpBranch && insn[14:12] == 3'b100;
  wire insn_bge = insn_opcode == OpBranch && insn[14:12] == 3'b101;
  wire insn_bltu = insn_opcode == OpBranch && insn[14:12] == 3'b110;
  wire insn_bgeu = insn_opcode == OpBranch && insn[14:12] == 3'b111;

  wire insn_lb = insn_opcode == OpLoad && insn[14:12] == 3'b000;
  wire insn_lh = insn_opcode == OpLoad && insn[14:12] == 3'b001;
  wire insn_lw = insn_opcode == OpLoad && insn[14:12] == 3'b010;
  wire insn_lbu = insn_opcode == OpLoad && insn[14:12] == 3'b100;
  wire insn_lhu = insn_opcode == OpLoad && insn[14:12] == 3'b101;

  wire insn_sb = insn_opcode == OpStore && insn[14:12] == 3'b000;
  wire insn_sh = insn_opcode == OpStore && insn[14:12] == 3'b001;
  wire insn_sw = insn_opcode == OpStore && insn[14:12] == 3'b010;

  wire insn_addi = insn_opcode == OpRegImm && insn[14:12] == 3'b000;
  wire insn_slti = insn_opcode == OpRegImm && insn[14:12] == 3'b010;
  wire insn_sltiu = insn_opcode == OpRegImm && insn[14:12] == 3'b011;
  wire insn_xori = insn_opcode == OpRegImm && insn[14:12] == 3'b100;
  wire insn_ori = insn_opcode == OpRegImm && insn[14:12] == 3'b110;
  wire insn_andi = insn_opcode == OpRegImm && insn[14:12] == 3'b111;

  wire insn_slli = insn_opcode == OpRegImm && insn[14:12] == 3'b001 && insn[31:25] == 7'd0;
  wire insn_srli = insn_opcode == OpRegImm && insn[14:12] == 3'b101 && insn[31:25] == 7'd0;
  wire insn_srai = insn_opcode == OpRegImm && insn[14:12] == 3'b101 && insn[31:25] == 7'b0100000;

  wire insn_add = insn_opcode == OpRegReg && insn[14:12] == 3'b000 && insn[31:25] == 7'd0;
  wire insn_sub  = insn_opcode == OpRegReg && insn[14:12] == 3'b000 && insn[31:25] == 7'b0100000;
  wire insn_sll = insn_opcode == OpRegReg && insn[14:12] == 3'b001 && insn[31:25] == 7'd0;
  wire insn_slt = insn_opcode == OpRegReg && insn[14:12] == 3'b010 && insn[31:25] == 7'd0;
  wire insn_sltu = insn_opcode == OpRegReg && insn[14:12] == 3'b011 && insn[31:25] == 7'd0;
  wire insn_xor = insn_opcode == OpRegReg && insn[14:12] == 3'b100 && insn[31:25] == 7'd0;
  wire insn_srl = insn_opcode == OpRegReg && insn[14:12] == 3'b101 && insn[31:25] == 7'd0;
  wire insn_sra  = insn_opcode == OpRegReg && insn[14:12] == 3'b101 && insn[31:25] == 7'b0100000;
  wire insn_or = insn_opcode == OpRegReg && insn[14:12] == 3'b110 && insn[31:25] == 7'd0;
  wire insn_and = insn_opcode == OpRegReg && insn[14:12] == 3'b111 && insn[31:25] == 7'd0;

  wire insn_mul    = insn_opcode == OpRegReg && insn[31:25] == 7'd1 && insn[14:12] == 3'b000;
  wire insn_mulh   = insn_opcode == OpRegReg && insn[31:25] == 7'd1 && insn[14:12] == 3'b001;
  wire insn_mulhsu = insn_opcode == OpRegReg && insn[31:25] == 7'd1 && insn[14:12] == 3'b010;
  wire insn_mulhu  = insn_opcode == OpRegReg && insn[31:25] == 7'd1 && insn[14:12] == 3'b011;
  wire insn_div    = insn_opcode == OpRegReg && insn[31:25] == 7'd1 && insn[14:12] == 3'b100;
  wire insn_divu   = insn_opcode == OpRegReg && insn[31:25] == 7'd1 && insn[14:12] == 3'b101;
  wire insn_rem    = insn_opcode == OpRegReg && insn[31:25] == 7'd1 && insn[14:12] == 3'b110;
  wire insn_remu   = insn_opcode == OpRegReg && insn[31:25] == 7'd1 && insn[14:12] == 3'b111;

  wire insn_ecall = insn_opcode == OpEnviron && insn[31:7] == 25'd0;
  wire insn_fence = insn_opcode == OpMiscMem;

  `include "RvDisassembler.sv"
  string disasm_string;
  always_comb begin
    disasm_string = rv_disasm(insn);
  end
  // HACK: get disasm_string to appear in GtkWave, which can apparently show only wire/logic...
  wire [(8*32)-1:0] disasm_wire;
  genvar i;
  for (i = 0; i < 32; i = i + 1) begin : gen_disasm
    assign disasm_wire[(((i+1))*8)-1:((i)*8)] = disasm_string[31-i];
  end

  // program counter
  logic [`REG_SIZE] pcNext, pcCurrent;
  always @(posedge clk) begin
    if (rst) begin
      pcCurrent <= 32'd0;
    end else begin
      pcCurrent <= pcNext;
    end
  end
  assign pc = pcCurrent;

  // cycle/insn counters
  logic [`REG_SIZE] cycles_current, num_insns_current;
  always @(posedge clk) begin
    if (rst) begin
      cycles_current <= 0;
      num_insns_current <= 0;
    end else begin
      cycles_current <= cycles_current + 1;
      if (!rst) begin
        num_insns_current <= num_insns_current + 1;
      end
    end
  end

  logic illegal_insn;

  always_comb begin
    illegal_insn = 1'b0;

    case (insn_opcode)
      OpLui: begin
        // TODO: start here by implementing lui
      end
      default: begin
        illegal_insn = 1'b1;
      end
    endcase
  end

endmodule

/**
  This memory module provides asynchronous reads. Writes are synchronous on the *negative* clock edge,
  so that they can take place within 1 processor clock cycle.
*/
module MemorySingleCycle #(
    parameter int NUM_WORDS = 512
) (
    input wire clk,
    input wire rst,

    // must always be aligned to a 4B boundary
    input wire [`REG_SIZE] addr0,

    // the value at memory location addr0
    output logic [`REG_SIZE] dout0,

    // must always be aligned to a 4B boundary
    input wire [`REG_SIZE] addr1,

    // the value at memory location addr1
    output logic [`REG_SIZE] dout1,

    // the value to be written to addr1, controlled by we1
    input wire [`REG_SIZE] din1,

    // Each bit determines whether to write the corresponding byte of din1 to memory location addr1.
    // E.g., 4'b1111 will write 4 bytes. 4'b0001 will write only the least-significant byte.
    input wire [3:0] we1
);

  // memory is arranged as an array of 4B words
  logic [`REG_SIZE] mem[NUM_WORDS];

  always_comb begin
    // memory addresses should always be 4B-aligned
    assert (addr0[1:0] == 2'b00);
    assert (addr1[1:0] == 2'b00);
  end

  localparam int AddrMsb = $clog2(NUM_WORDS) + 1;
  localparam int AddrLsb = 2;

  assign dout0 = mem[{addr0[AddrMsb:AddrLsb]}];
  assign dout1 = mem[{addr1[AddrMsb:AddrLsb]}];

  always @(negedge clk) begin
    if (rst) begin
    end else begin
      if (we1[0]) begin
        mem[addr1[AddrMsb:AddrLsb]][7:0] = din1[7:0];
      end
      if (we1[1]) begin
        mem[addr1[AddrMsb:AddrLsb]][15:8] = din1[15:8];
      end
      if (we1[2]) begin
        mem[addr1[AddrMsb:AddrLsb]][23:16] = din1[23:16];
      end
      if (we1[3]) begin
        mem[addr1[AddrMsb:AddrLsb]][31:24] = din1[31:24];
      end
    end
  end
endmodule

module RiscvProcessor (
    input  wire  clk,
    input  wire  rst,
    output logic halt
);

  wire [`REG_SIZE] pc, insn, mem_data_addr, mem_data_loaded_value, mem_data_to_write;
  wire [3:0] mem_data_we;

  MemorySingleCycle #(
      .NUM_WORDS(16384)
  ) mem (
      .clk  (clk),
      .rst  (rst),
      // addr0 is a read-only port
      .addr0(pc),
      .dout0(insn),
      // addr1 is a read-write port
      .addr1(mem_data_addr),
      .dout1(mem_data_loaded_value),
      .din1 (mem_data_to_write),
      .we1  (mem_data_we)
  );

  DatapathSingleCycle datapath (
      .clk(clk),
      .rst(rst),
      .pc(pc),
      .insn(insn),
      .addr1(mem_data_addr),
      .dout1(mem_data_loaded_value),
      .din1(mem_data_to_write),
      .we1(mem_data_we),
      .halt(halt)
  );

endmodule
