`default_nettype none
`timescale 1ns / 1ps

// registers are 32 bits in RV32
`define REG_SIZE 31:0

// insns are 32 bits in RV32IM
`define INSN_SIZE 31:0

`define RESP_OK 2'b00


`ifdef SYNTHESIS
`include "MyClockGen.v"
`endif

`include "DatapathPipelinedCache.sv"
`include "system/hdmi/hdmi_video.v"
`include "system/hdmi/vga_video.v"
`include "system/hdmi/vga2dvid.v"
`include "system/hdmi/fake_differential.v"
`include "system/hdmi/tmds_encoder.v"
`include "system/usb/usb_hid_host.v"
`include "../hw3-singlecycle/system/debouncer.v"

// FULL_SIZE_MEM means 32KB memory, FULL_SIZE_DISPLAY means 320x240 frame buffer
// non-FULL_SIZE means 4KB memory and 40x30 frame buffer, respectively
`define FULL_SIZE_MEM
`define FULL_SIZE_DISPLAY

module SystemResourceCheck (
    input wire external_clk_25MHz,
    input wire [6:0] btn,
    output wire [7:0] led
);

wire clk, clk_locked;
MyClockGen clock_gen (
  .input_clk_25MHz(external_clk_25MHz),
  .clk_proc(clk),
  .locked(clk_locked)
);
wire rst = !clk_locked;

axi_if axi_data_cache ();
// memory is dual-ported, to connect to both datapath and D$
axi_if axi_mem_ro ();
axi_if axi_mem_rw ();

AxilMemory #(.NUM_WORDS(8192)) memory (
  .ACLK(clk),
  .ARESETn(~rst),
  .port_ro(axi_mem_ro.subord),
  .port_rw(axi_mem_rw.subord)
);

  AxilCache #(
    .BLOCK_SIZE_BITS(32),
    .NUM_SETS(16)) dcache (
    .ACLK(clk),
    .ARESETn(~rst),
    .proc(axi_data_cache.subord),
    .mem(axi_mem_rw.manager)
  );

  DatapathPipelinedCache datapath (
      .clk(clk),
      .rst(rst),
      .icache(axi_mem_ro.manager),
      .dcache(axi_data_cache.manager),
      .halt(led[0])
  );
endmodule

/** NB: this module was generated by ecppll, do not edit manually */
module DemoClockGen
(
    input input_clk_25MHz, // 25 MHz, 0 deg
    output clk_125MHz, // 125 MHz, 0 deg
    output clk_25MHz, // 25 MHz, 0 deg
    output clk_12MHz, // 12.0192 MHz, 0 deg
    output locked
);
wire clkfb;
(* FREQUENCY_PIN_CLKI="25" *)
(* FREQUENCY_PIN_CLKOP="125" *)
(* FREQUENCY_PIN_CLKOS="25" *)
(* FREQUENCY_PIN_CLKOS2="12.0192" *)
(* ICP_CURRENT="12" *) (* LPF_RESISTOR="8" *) (* MFG_ENABLE_FILTEROPAMP="1" *) (* MFG_GMCREF_SEL="2" *)
EHXPLLL #(
        .PLLRST_ENA("DISABLED"),
        .INTFB_WAKE("DISABLED"),
        .STDBY_ENABLE("DISABLED"),
        .DPHASE_SOURCE("DISABLED"),
        .OUTDIVIDER_MUXA("DIVA"),
        .OUTDIVIDER_MUXB("DIVB"),
        .OUTDIVIDER_MUXC("DIVC"),
        .OUTDIVIDER_MUXD("DIVD"),
        .CLKI_DIV(1),
        .CLKOP_ENABLE("ENABLED"),
        .CLKOP_DIV(5),
        .CLKOP_CPHASE(2),
        .CLKOP_FPHASE(0),
        .CLKOS_ENABLE("ENABLED"),
        .CLKOS_DIV(25),
        .CLKOS_CPHASE(2),
        .CLKOS_FPHASE(0),
        .CLKOS2_ENABLE("ENABLED"),
        .CLKOS2_DIV(52),
        .CLKOS2_CPHASE(2),
        .CLKOS2_FPHASE(0),
        .FEEDBK_PATH("INT_OP"),
        .CLKFB_DIV(5)
    ) pll_i (
        .RST(1'b0),
        .STDBY(1'b0),
        .CLKI(input_clk_25MHz),
        .CLKOP(clk_125MHz),
        .CLKOS(clk_25MHz),
        .CLKOS2(clk_12MHz),
        .CLKFB(clkfb),
        .CLKINTFB(clkfb),
        .PHASESEL0(1'b0),
        .PHASESEL1(1'b0),
        .PHASEDIR(1'b1),
        .PHASESTEP(1'b1),
        .PHASELOADREG(1'b1),
        .PLLWAKESYNC(1'b0),
        .ENCLKOP(1'b0),
        .LOCK(locked)
	);
endmodule

module MemoryMap (
    input wire ACLK,
    input wire ARESETn,
    axi_if.subord proc,
    axi_if.manager cache,
    input wire clk_25MHz,
    input wire clk_125MHz,
    input wire clk_12MHz,
    input wire clk_locked,
    input wire [6:0] btn,
    output wire [7:0] led,
    output wire [3:0] gpdi_dp,
    output wire [3:0] gpdi_dn,
    inout wire usb_fpga_bd_dn,
    inout wire usb_fpga_bd_dp
);

  // This module is a "bump on the wire", a (conceptually) combinational circuit between proc and cache.

  localparam int MmapButtons   = 32'hFF00_1000;
  localparam int MmapLeds      = 32'hFF00_2000;
  //localparam int MmapUartRead    = 32'hFF00_3000;
  //localparam int MmapUartWrite    = 32'hFF00_3001;
  localparam int MmapUsb       = 32'hFF00_4000;
  localparam int MmapRng       = 32'hFF00_5000;
  localparam int MmapHdmiStart = 32'hFF10_0000;
  `ifdef FULL_SIZE_DISPLAY
  localparam bit[9:0] HdmiWidth = 320;
  localparam bit[9:0] HdmiHeight = 240;
  `else
  localparam bit[9:0] HdmiWidth = 40;
  localparam bit[9:0] HdmiHeight = 30;
  `endif
  localparam int HdmiPixels = HdmiHeight * HdmiWidth;
  localparam int HdmiPixelSizeBits = 8;
  localparam bit[9:0] HdmiFrameBufferScale = 640 / HdmiWidth;
  localparam int HdmiFrameBufferScaleShift = $clog2(HdmiFrameBufferScale);
  localparam int MmapHdmiEnd = MmapHdmiStart + (HdmiPixels * (HdmiPixelSizeBits / 8));

  localparam bit True = 1'b1;
  localparam bit False = 1'b0;

  assign cache.ARADDR = proc.ARADDR;
  assign cache.ARVALID = is_read ? False : proc.ARVALID;  // hide request from the cache
  assign cache.ARPROT = proc.ARPROT;
  assign proc.ARREADY = cache.ARREADY;
  assign cache.RREADY = proc.RREADY;
  assign proc.RVALID = was_read ? True : cache.RVALID;
  assign proc.RDATA =
    was_board_button ? {{proc.ADDR_WIDTH - 7{1'b0}}, btn} :
    was_usb ? {{proc.DATA_WIDTH - 10{1'b0}}, usb_buttons} :
    was_rng ? rng_state : cache.RDATA;
  assign proc.RRESP = cache.RRESP;

  assign cache.AWADDR = proc.AWADDR;

  assign cache.AWVALID = is_write ? False : proc.AWVALID;  // hide request from the cache
  assign cache.WVALID = is_write ? False : proc.WVALID;
  assign proc.AWREADY = cache.AWREADY;
  assign cache.AWPROT = proc.AWPROT;
  assign cache.WDATA = proc.WDATA;
  assign cache.WSTRB = proc.WSTRB;
  assign proc.WREADY = cache.WREADY;
  assign cache.BREADY = proc.BREADY;
  assign proc.BVALID = was_write ? True : cache.BVALID;
  assign proc.BRESP = cache.BRESP;

  logic [proc.ADDR_WIDTH-1:0] last_araddr, last_awaddr;
  logic [proc.DATA_WIDTH-1:0] last_wdata;
  logic [(proc.DATA_WIDTH/8)-1:0] last_wstrb;
  logic last_arvalid, last_arready, last_awvalid, last_awready, last_wvalid, last_wready;

  wire is_axi_read = proc.ARVALID && cache.ARREADY;
  wire is_board_button = is_axi_read && (proc.ARADDR == MmapButtons);
  wire is_usb = is_axi_read && (proc.ARADDR == MmapUsb);
  wire is_rng = is_axi_read && (proc.ARADDR == MmapRng);
  wire is_read = is_board_button || is_usb || is_rng;
  wire was_axi_read = last_arvalid && last_arready;
  wire was_board_button = was_axi_read && (last_araddr == MmapButtons);
  wire was_usb = was_axi_read && (last_araddr == MmapUsb);
  wire was_rng = was_axi_read && (last_araddr == MmapRng);
  wire was_read = was_board_button || was_usb || was_rng;

  wire is_axi_write = proc.AWVALID && cache.AWREADY && proc.WVALID && cache.WREADY;
  wire is_led = is_axi_write && (proc.AWADDR == MmapLeds);
  wire is_hdmi = is_axi_write && (MmapHdmiStart <= proc.AWADDR && proc.AWADDR < MmapHdmiEnd);
  wire is_write = is_led || is_hdmi;
  wire was_axi_write = last_awvalid && last_awready && last_wvalid && last_wready;
  wire was_led = was_axi_write && (last_awaddr == MmapLeds);
  wire was_hdmi = was_axi_write && (MmapHdmiStart <= last_awaddr && last_awaddr < MmapHdmiEnd);
  wire was_write = was_led || was_hdmi;

  always_ff @(posedge ACLK) begin
    if (!ARESETn) begin
      last_araddr  <= 0;
      last_arvalid <= False;
      last_arready <= False;

      last_awaddr  <= 0;
      last_awvalid <= False;
      last_awready <= False;
      last_wdata   <= 0;
      last_wstrb   <= 0;
      last_wvalid  <= False;
      last_wready <= False;
    end else begin
      last_araddr  <= proc.ARADDR;
      last_arvalid <= proc.ARVALID;
      last_arready <= cache.ARREADY;

      last_awaddr  <= proc.AWADDR;
      last_awvalid <= proc.AWVALID;
      last_awready <= cache.AWREADY;
      last_wdata   <= proc.WDATA;
      last_wstrb   <= proc.WSTRB;
      last_wvalid  <= proc.WVALID;
      last_wready  <= cache.WREADY;
    end
  end

  // NB: Buttons are implemented above as mux on RDATA

  // Random Number Generator: a linear-feedback shift register

  logic [31:0] rng_state;
  logic feedback;
  always_ff @(posedge ACLK) begin
    if (!ARESETn) begin
      rng_state <= 12345;
    end else begin
      feedback <= rng_state[0] ^ rng_state[1] ^ rng_state[21] ^ rng_state[31]; // XOR taps
      rng_state <= {rng_state[30:0], feedback}; // Shift left and insert feedback
    end
  end

  // LEDs

  logic [7:0] led_state;
  assign led = led_state[7:0];
  always_ff @(posedge ACLK) begin
    if (!ARESETn) begin
      led_state <= 0;
    end else begin
      if (was_led) begin
        led_state <= last_wdata[7:0];
      end
    end
  end

  // USB

  wire [1:0] usb_type;
  wire [7:0] key_modifiers, key1, key2, key3, key4;
  wire [7:0] mouse_btn;
  wire signed [7:0] mouse_dx, mouse_dy;
  wire [63:0] hid_report;
  wire usb_report, usb_conerr;
  wire game_l, game_r, game_u, game_d, game_a, game_b, game_x, game_y;
  wire game_select, game_start;
  wire [9:0] usb_buttons = {
    game_l, game_r, game_u, game_d, game_a, game_b, game_x, game_y, game_select, game_start
  };

`ifdef SYNTHESIS
  usb_hid_host usb (
      .usbclk(clk_12MHz),
      .usbrst_n(ARESETn),
      .usb_dm(usb_fpga_bd_dn),
      .usb_dp(usb_fpga_bd_dp),
      .typ(usb_type),
      .report(usb_report),
      .key_modifiers(key_modifiers),
      .key1(key1),
      .key2(key2),
      .key3(key3),
      .key4(key4),
      .mouse_btn(mouse_btn),
      .mouse_dx(mouse_dx),
      .mouse_dy(mouse_dy),
      .game_l(game_l),
      .game_r(game_r),
      .game_u(game_u),
      .game_d(game_d),
      .game_a(game_a),
      .game_b(game_b),
      .game_x(game_x),
      .game_y(game_y),
      .game_sel(game_select),
      .game_sta(game_start),
      .conerr(usb_conerr),
      .dbg_hid_report(hid_report)
  );
`endif

  // HDMI frame buffer

//   localparam bit [7:0] Black = 8'b000_000_00;
//   localparam bit [7:0] Red   = 8'b111_000_00;
  localparam bit [7:0] White = 8'b111_111_11;
//   localparam bit [7:0] Teal  = 8'b000_111_10;

  logic [HdmiPixelSizeBits-1:0] frame_buffer[HdmiWidth * HdmiHeight];
  initial begin
    for (integer i = 0; i < HdmiPixels; i = i + 1) begin
        frame_buffer[i] = White;
    end
  end
  always_ff @(posedge ACLK) begin
    if (ARESETn) begin
      if (was_hdmi) begin
        case (last_wstrb)
        4'b0001: begin
            frame_buffer[last_awaddr-MmapHdmiStart] <= last_wdata[7:0];
        end
        4'b0010: begin
            frame_buffer[(last_awaddr-MmapHdmiStart)+1] <= last_wdata[15:8];
        end
        4'b0100: begin
            frame_buffer[(last_awaddr-MmapHdmiStart)+2] <= last_wdata[23:16];
        end
        4'b1000: begin
            frame_buffer[(last_awaddr-MmapHdmiStart)+3] <= last_wdata[31:24];
        end
        default: begin end
        endcase
      end
    end
  end

  wire [9:0] raw_x, raw_y, raw_x_scaled, raw_y_scaled;
  assign raw_x_scaled = raw_x >> HdmiFrameBufferScaleShift[3:0];
  assign raw_y_scaled = raw_y >> HdmiFrameBufferScaleShift[3:0];
  wire [9:0] x = raw_x_scaled < HdmiWidth ? raw_x_scaled : HdmiWidth - 1;
  wire [8:0] y = raw_y_scaled < HdmiHeight ? raw_y_scaled[8:0] : 9'd119;

`ifdef FULL_SIZE_DISPLAY
  // NB: use this for 320x240 display
  wire [16:0] fb_index = ({8'd0, y} * {7'd0, HdmiWidth}) + {7'd0, x};
`else
  // NB: use this for 40x30 display
  wire [10:0] fb_index = ({2'd0, y} * {1'd0, HdmiWidth}) + {1'd0, x};
`endif

  logic [HdmiPixelSizeBits-1:0] color8;
  always_ff @(posedge clk_25MHz) begin
    if (!ARESETn) begin
      color8 <= 0;
    end else begin
      color8 <= frame_buffer[fb_index];
    end
  end

  // scale from 8-bit color to 24-bit color
  wire [7:0] red24   = {color8[7:5], color8[7:5], color8[7:6]};
  wire [7:0] green24 = {color8[4:2], color8[4:2], color8[4:3]};
  wire [7:0] blue24  = {color8[1:0], color8[1:0], color8[1:0], color8[1:0]};

  wire [23:0] color24 = {red24, green24, blue24};
`ifdef SYNTHESIS
  hdmi_video hdmi_video (
      .clk_25MHz(clk_25MHz),
      .clk_125MHz(clk_125MHz),
      .clk_locked(clk_locked),
      .x(raw_x),
      .y(raw_y),
      .color(color24),
      .gpdi_dp(gpdi_dp),
      .gpdi_dn(gpdi_dn)
  );
`endif

endmodule

module SystemDemo (
    input wire external_clk_25MHz,
    input wire [6:0] btn,
    output wire [7:0] led,
    output wire [3:0] gpdi_dp,
    output wire [3:0] gpdi_dn,
    inout wire  usb_fpga_bd_dn,
    inout wire  usb_fpga_bd_dp,
    output wire ftdi_rxd, // from FPGA to host
    inout wire gpdi_sda,
    output wire gpdi_scl
);

  // NB: btn[0] is active-low: it sends 1 when not pressed, and 0 when pressed
  wire rst_n;
`ifdef SYNTHESIS
  wire [30:0] ignore;
  debouncer #(.NIN(1)) db (
      .i_clk(clk_proc),
      .i_in(btn[0]),
      .o_debounced(rst_n),
      .o_debug(ignore)
  );
`else
  assign rst_n = btn[0];
`endif

  localparam bit True = 1'b1;
//   localparam bit False = 1'b0;
  wire clk_25MHz, clk_125MHz, clk_12MHz, clk_proc, clk_locked, demo_clocks_locked;

`ifdef SYNTHESIS
  MyClockGen clock_gen (
    .input_clk_25MHz(external_clk_25MHz),
    .clk_proc(clk_proc),
    .locked(clk_locked)
    );

    DemoClockGen demo_clock_gen (
    .input_clk_25MHz(external_clk_25MHz),
    .locked(demo_clocks_locked),
    .clk_125MHz(clk_125MHz),
    .clk_25MHz(clk_25MHz),
    .clk_12MHz(clk_12MHz)
);
`else
    assign clk_25MHz  = external_clk_25MHz;
    assign clk_proc   = external_clk_25MHz;
    assign clk_125MHz = external_clk_25MHz;
    assign clk_locked = True;
`endif
  wire rst = !rst_n || !clk_locked || !demo_clocks_locked;

  axi_if axi_data_cache ();
  axi_if axi_data_mmap ();
  axi_if axi_insn_cache ();
  // memory is dual-ported, to connect to both I$ and D$
  axi_if axi_mem_a ();
  axi_if axi_mem_b ();

`ifdef FULL_SIZE_MEM
  AxilMemory #(.NUM_WORDS(8192)) the_mem
`else
  AxilMemory #(.NUM_WORDS(2048)) the_mem
`endif
  (
      .ACLK(clk_proc),
      .ARESETn(~rst),
      .port_ro(axi_mem_a.subord),
      .port_rw(axi_mem_b.subord)
  );

  MemoryMap mmap (
      .ACLK(clk_proc),
      .ARESETn(~rst),
      .proc(axi_data_mmap.subord),
      .cache(axi_data_cache.manager),
      .clk_25MHz(clk_25MHz),
      .clk_125MHz(clk_125MHz),
      .clk_locked(clk_locked),
      .btn(btn),
      .led(led),
      .gpdi_dp(gpdi_dp),
      .gpdi_dn(gpdi_dn),
      .usb_fpga_bd_dn(usb_fpga_bd_dn),
      .usb_fpga_bd_dp(usb_fpga_bd_dp)
  );

  AxilCache #(
      .BLOCK_SIZE_BITS(32),
      .NUM_SETS(64)
  ) dcache (
      .ACLK(clk_proc),
      .ARESETn(~rst),
      .proc(axi_data_cache.subord),
      .mem(axi_mem_b.manager)
  );

  wire halt;

  DatapathPipelinedCache datapath (
      .clk(clk_proc),
      .rst(rst),
      .icache(axi_mem_a.manager),
      .dcache(axi_data_mmap.manager),
      .halt(halt)
  );

endmodule

module SystemSim (
    input wire external_clk_25MHz,
    input wire rst,
    input wire [6:0] btn,
    output wire [7:0] led,
    output wire [3:0] gpdi_dp,
    output wire [3:0] gpdi_dn,
    inout wire  usb_fpga_bd_dn,
    inout wire  usb_fpga_bd_dp,
    output wire ftdi_rxd // from FPGA to host
);

  localparam bit True = 1'b1;
//   localparam bit False = 1'b0;
  wire clk_25MHz, clk_125MHz, clk_proc, clk_locked;

  assign clk_25MHz  = external_clk_25MHz;
  assign clk_proc   = external_clk_25MHz;
  assign clk_125MHz = external_clk_25MHz;
  assign clk_locked = True;

  axi_if axi_data_cache ();
  axi_if axi_data_mmap ();
  axi_if axi_insn_cache ();
  // memory is dual-ported, to connect to both I$ and D$
  axi_if axi_mem_a ();
  axi_if axi_mem_b ();

  wire [7:0] fake_led, fake_led2;

`ifdef FULL_SIZE_MEM
  AxilMemory #(.NUM_WORDS(8192)) the_mem
`else
  AxilMemory #(.NUM_WORDS(2048)) the_mem
`endif
  (
      .ACLK(clk_proc),
      .ARESETn(~rst),
      .port_ro(axi_mem_a.subord),
      .port_rw(axi_mem_b.subord)
  );

  MemoryMap mmap (
      .ACLK(clk_proc),
      .ARESETn(~rst),
      .proc(axi_data_mmap.subord),
      .cache(axi_data_cache.manager),
      .clk_25MHz(clk_25MHz),
      .clk_125MHz(clk_125MHz),
      .clk_locked(clk_locked),
      .btn(btn),
      .led(fake_led),
      .gpdi_dp(gpdi_dp),
      .gpdi_dn(gpdi_dn),
      .usb_fpga_bd_dn(usb_fpga_bd_dn),
      .usb_fpga_bd_dp(usb_fpga_bd_dp)
  );

  AxilCache #(
      .BLOCK_SIZE_BITS(32),
      .NUM_SETS(16)
  ) icache (
      .ACLK(clk_proc),
      .ARESETn(~rst),
      .proc(axi_insn_cache.subord),
      .mem(axi_mem_a.manager)
  );

  AxilCache #(
      .BLOCK_SIZE_BITS(32),
      .NUM_SETS(16)
  ) dcache (
      .ACLK(clk_proc),
      .ARESETn(~rst),
      .proc(axi_data_cache.subord),
      .mem(axi_mem_b.manager)
  );

  wire halt;
  wire [`REG_SIZE] trace_writeback_pc;
  wire [`INSN_SIZE] trace_writeback_insn;
  wire cycle_status_e trace_writeback_cycle_status;

  // localparam int MmapButtons   = 32'hFF00_1000;
  localparam int MmapLeds      = 32'hFF00_2000;
  //localparam int MmapUartRead    = 32'hFF00_3000;
  //localparam int MmapUartWrite    = 32'hFF00_3001;
  // localparam int MmapUsb       = 32'hFF00_4000;
  // localparam int MmapRng       = 32'hFF00_5000;
  localparam int MmapHdmiStart = 32'hFF10_0000;
  `ifdef FULL_SIZE_DISPLAY
  localparam bit[9:0] HdmiWidth = 320;
  localparam bit[9:0] HdmiHeight = 240;
  `else
  localparam bit[9:0] HdmiWidth = 40;
  localparam bit[9:0] HdmiHeight = 30;
  `endif
  localparam int HdmiPixels = HdmiHeight * HdmiWidth;
  localparam int HdmiPixelSizeBits = 8;
  // localparam bit[9:0] HdmiFrameBufferScale = 640 / HdmiWidth;
  // localparam int HdmiFrameBufferScaleShift = $clog2(HdmiFrameBufferScale);
  localparam int MmapHdmiEnd = MmapHdmiStart + (HdmiPixels * (HdmiPixelSizeBits / 8));

  wire is_write_to_read_only = axi_data_cache.manager.AWVALID &&
        axi_data_cache.manager.AWADDR[14:0] <= 15'h6000 &&
        axi_data_cache.manager.AWADDR != MmapLeds &&
        (axi_data_cache.manager.AWADDR < MmapHdmiStart || axi_data_cache.manager.AWADDR > MmapHdmiEnd);

  DatapathPipelinedCache datapath (
      .clk(clk_proc),
      .rst(rst),
      .icache(axi_insn_cache.manager),
      .dcache(axi_data_mmap.manager),
      // .dcache(axi_data_cache.manager),
      .halt(halt),
      .trace_writeback_pc(trace_writeback_pc),
      .trace_writeback_insn(trace_writeback_insn),
      .trace_writeback_cycle_status(trace_writeback_cycle_status)
  );

endmodule
