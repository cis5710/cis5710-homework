/**
 * This enum is used to classify the work happening in each cycle, to validate
 * datapath timing. For single-cycle designs, the datapath never stalls. With
 * multi-cycle designs, the possibility of stall cycles arises. For pipelined
 * designs, we classify only the work happening in the Writeback stage,
 * identifying if a valid insn is present or, if it is a stall cycle instead,
 * the reason for the stall. These values are compared against the trace-*.json
 * files to ensure that the datapath is doing the correct operation in each
 * cycle.
 *
 * For pipelined designs, you will need to set these values at various places
 * within your pipeline, and propagate them through the stages until they reach
 * Writeback where they can be checked. Note that MULTIPLE stall conditions may
 * be present in a single cycle. All relevant stall conditions should be ORed
 * together.
 */
typedef enum {
  /** invalid value, this should never appear after the initial reset sequence completes */
  CYCLE_INVALID = 0,
  /** not a stall cycle, a valid insn is in Writeback */
  CYCLE_NO_STALL = 1,

  // the values below are only needed in HW4 and later
              
  /** a stall cycle that arose from waiting for a multi-cycle div/rem insn */
  CYCLE_DIV = 2,

  // the values below are only needed in HW5A and later
              
  /** a stall cycle that arose from the pipeline being initially empty */
  CYCLE_RESET = 4,
  /** a stall cycle that arose from a taken branch/jump */
  CYCLE_TAKEN_BRANCH = 8,

  // the values below are only needed in HW5B and later

  /** a stall cycle that arose from a load-to-use stall */
  CYCLE_LOAD2USE = 16,
  /** NOT CURRENTLY USED */
  CYCLE_DIV2USE = 32,
  /** NOT CURRENTLY USED: a stall cycle that arose from a fence.i insn */
  CYCLE_FENCEI = 64,

  // the values below are only needed in HW6B

  /** a stall cycle that arose from an insn cache miss */
  CYCLE_ICACHE_MISS = 128,
  /** a stall cycle that arose from a data cache miss */
  CYCLE_DCACHE_MISS = 256

} cycle_status_e;
